//
// Copyright (c) 2016, Intel Corporation
// All rights reserved.
//
// Redistribution and use in source and binary forms, with or without
// modification, are permitted provided that the following conditions are met:
//
// Redistributions of source code must retain the above copyright notice, this
// list of conditions and the following disclaimer.
//
// Redistributions in binary form must reproduce the above copyright notice,
// this list of conditions and the following disclaimer in the documentation
// and/or other materials provided with the distribution.
//
// Neither the name of the Intel Corporation nor the names of its contributors
// may be used to endorse or promote products derived from this software
// without specific prior written permission.
//
// THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS"
// AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE
// IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE
// ARE DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT OWNER OR CONTRIBUTORS BE
// LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR
// CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF
// SUBSTITUTE GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS
// INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN
// CONTRACT, STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
// ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE
// POSSIBILITY OF SUCH DAMAGE.

//
// test_random configuration.  These are in ifdefs so they can be overridden
// by command line definitions.
//

`ifndef MPF_CONF_SORT_READ_RESPONSES
  `define MPF_CONF_SORT_READ_RESPONSES 1
`endif

`ifndef MPF_CONF_PRESERVE_WRITE_MDATA
  `define MPF_CONF_PRESERVE_WRITE_MDATA 1
`endif

`ifndef MPF_CONF_ENABLE_VTP
  `define MPF_CONF_ENABLE_VTP 1
`endif

// Software translation service
//`define MPF_CONF_VTP_PT_MODE_SOFTWARE_SERVICE

`ifndef MPF_CONF_ENABLE_VC_MAP
  `define MPF_CONF_ENABLE_VC_MAP 1
`endif

`ifndef MPF_CONF_ENFORCE_WR_ORDER
  `define MPF_CONF_ENFORCE_WR_ORDER 1
`endif

`ifndef MPF_CONF_ENABLE_PARTIAL_WRITES
  `define MPF_CONF_ENABLE_PARTIAL_WRITES 1
`endif
`ifndef MPF_CONF_PARTIAL_WRITE_MODE
  `define MPF_CONF_PARTIAL_WRITE_MODE "BYTE_RANGE"
`endif
