//
// MPF's view of CCI expressed as a SystemVerilog interface.
//

`ifndef CCI_MPF_IF_VH
`define CCI_MPF_IF_VH

`include "cci_mpf_platform.vh"

import cci_mpf_if_pkg::*;
import ccip_if_funcs_pkg::*;

`endif //  CCI_MPF_IF_VH
