// lpbk1_RdRspRAM2PORT.v

// Generated using ACDS version 15.1 192

`timescale 1 ps / 1 ps
module lpbk1_RdRspRAM2PORT (
		input  wire [533:0] data,      //  ram_input.datain
		input  wire [8:0]   wraddress, //           .wraddress
		input  wire [8:0]   rdaddress, //           .rdaddress
		input  wire         wren,      //           .wren
		input  wire         clock,     //           .clock
		output wire [533:0] q          // ram_output.dataout
	);

	lpbk1_RdRspRAM2PORT_ram_2port_151_davj2sq ram_2port_0 (
		.data      (data),      //  ram_input.datain
		.wraddress (wraddress), //           .wraddress
		.rdaddress (rdaddress), //           .rdaddress
		.wren      (wren),      //           .wren
		.clock     (clock),     //           .clock
		.q         (q)          // ram_output.dataout
	);

endmodule
