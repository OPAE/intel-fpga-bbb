// feeder_ram_512_256.v

// Generated using ACDS version 15.1 185

`timescale 1 ps / 1 ps
module feeder_ram_512_256 # (
	SIZE = 512
	) (
		input  wire [511:0]              data,      //  ram_input.datain
		input  wire [$clog2(SIZE)-1:0]   wraddress, //           .wraddress
		input  wire [$clog2(SIZE*2)-1:0] rdaddress, //           .rdaddress
		input  wire                      wren,      //           .wren
		input  wire                      clock,     //           .clock
		input  wire                      rden,      //           .rden
		output wire [255:0]              q          // ram_output.dataout
	);

	feeder_ram_512_256_ram_2port_151_i4icjwq # (SIZE) ram_2port_0 (
		.data      (data),      //  ram_input.datain
		.wraddress (wraddress), //           .wraddress
		.rdaddress (rdaddress), //           .rdaddress
		.wren      (wren),      //           .wren
		.clock     (clock),     //           .clock
		.rden      (rden),      //           .rden
		.q         (q)          // ram_output.dataout
	);

endmodule
