//
// Copyright (c) 2020, Intel Corporation
// All rights reserved.
//
// Redistribution and use in source and binary forms, with or without
// modification, are permitted provided that the following conditions are met:
//
// Redistributions of source code must retain the above copyright notice, this
// list of conditions and the following disclaimer.
//
// Redistributions in binary form must reproduce the above copyright notice,
// this list of conditions and the following disclaimer in the documentation
// and/or other materials provided with the distribution.
//
// Neither the name of the Intel Corporation nor the names of its contributors
// may be used to endorse or promote products derived from this software
// without specific prior written permission.
//
// THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS"
// AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE
// IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE
// ARE DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT OWNER OR CONTRIBUTORS BE
// LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR
// CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF
// SUBSTITUTE GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS
// INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN
// CONTRACT, STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
// ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE
// POSSIBILITY OF SUCH DAMAGE.

//
// Translate addresses for a single DMA request channel.
//

`include "cci_mpf_if.vh"

module mpf_vtp_translate_chan
  #(
    // Return results in request order if non-zero
    parameter ORDERED = 1,

    // Requests pass through the module as opaque values. Set the size
    // to match the opaque_* ports.
    parameter N_OPAQUE_BITS = 0
    )
   (
    input  logic clk,
    input  logic reset,

    output logic rsp_valid,
    output logic [N_OPAQUE_BITS-1 : 0] opaque_rsp,
    input  logic deq_en,

    // New request is accepted when req_valid and not full. req_valid is
    // ignored when VTP is full.
    input  logic req_valid,
    input  logic [N_OPAQUE_BITS-1 : 0] opaque_req,
    output logic full,

    // Request: commands to VTP (e.g. address to translate)
    input  mpf_vtp_pkg::t_mpf_vtp_port_wrapper_req vtp_req,
    // Response from VTP (e.g. whether translation was successful)
    output mpf_vtp_pkg::t_mpf_vtp_port_wrapper_rsp vtp_rsp,
    mpf_vtp_port_if.to_slave vtp_port
    );

    import mpf_vtp_pkg::*;

    logic vtp_notFull;
    assign full = ~vtp_notFull;

    t_mpf_vtp_req_tag vtp_reqIdx;
    t_mpf_vtp_req_tag vtp_rspIdx;

    // VTP assigns the request a unique ID while in flight (reqIdx). The
    // ID will be returned with the response (rspIdx), making it easy to
    // manage storage of request opaque data.
    generate
        if (ORDERED != 0)
        begin : o
            mpf_svc_vtp_port_wrapper_ordered
              tr
               (
                .clk,
                .reset,

                .vtp_port,
                .reqEn(req_valid && vtp_notFull),
                .req(vtp_req),
                .notFull(vtp_notFull),
                .reqIdx(vtp_reqIdx),

                .rspValid(rsp_valid),
                .rsp(vtp_rsp),
                .rspDeqEn(deq_en),
                .rspIdx(vtp_rspIdx)
                );
        end
        else
        begin : u
            mpf_svc_vtp_port_wrapper_unordered
              tr
               (
                .clk,
                .reset,

                .vtp_port,
                .reqEn(req_valid && vtp_notFull),
                .req(vtp_req),
                .notFull(vtp_notFull),
                .reqIdx(vtp_reqIdx),

                .rspValid(rsp_valid),
                .rsp(vtp_rsp),
                .rspDeqEn(deq_en),
                .rspIdx(vtp_rspIdx)
                );
        end
    endgenerate

    // Hold the opaque request during lookup. The VTP port wrapper provides
    // up to MPF_VTP_MAX_SVC_REQS indices. The addresses used for storage are
    // generated by the VTP port as part of its request tracking logic.
    cci_mpf_prim_lutram
      #(
        .N_ENTRIES(MPF_VTP_MAX_SVC_REQS),
        .N_DATA_BITS(N_OPAQUE_BITS)
        )
      tr_meta
       (
        .clk,
        .reset,

        .raddr(vtp_rspIdx),
        .rdata(opaque_rsp),

        .wen(req_valid && vtp_notFull),
        .waddr(vtp_reqIdx),
        .wdata(opaque_req)
        );


    //
    // Debugging
    //

    // synthesis translate_off
    always_ff @(posedge clk)
    begin
        if (! reset)
        begin
            if (deq_en && vtp_rsp.error)
            begin
                $display("%m VTP: %0t Translation error from VA 0x%x",
                         $time,
                         {vtp_rsp.addr, 6'b0});
            end
        end
    end
    // synthesis translate_on

endmodule // mpf_vtp_translate_chan_ordered
