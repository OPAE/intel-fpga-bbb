// dot16_result_fifo.v

// Generated using ACDS version 15.1 193

`timescale 1 ps / 1 ps
module dot16_result_fifo #(
  DATA_WIDTH = 32
) (
		input  wire [DATA_WIDTH-1:0]  data,        //  fifo_input.datain
		input  wire                   wrreq,       //            .wrreq
		input  wire                   rdreq,       //            .rdreq
		input  wire                   clock,       //            .clk
		input  wire                   sclr,        //            .sclr
		output wire [DATA_WIDTH-1:0]  q,           // fifo_output.dataout
		output wire [9:0]             usedw,       //            .usedw
		output wire                   full,        //            .full
		output wire                   empty,       //            .empty
		output wire                   almost_full  //            .almost_full
	);

	dot16_result_fifo_fifo_151_myzccvq # (
    .DATA_WIDTH (DATA_WIDTH)
  ) fifo_0 (
		.data        (data),        //  fifo_input.datain
		.wrreq       (wrreq),       //            .wrreq
		.rdreq       (rdreq),       //            .rdreq
		.clock       (clock),       //            .clk
		.sclr        (sclr),        //            .sclr
		.q           (q),           // fifo_output.dataout
		.usedw       (usedw),       //            .usedw
		.full        (full),        //            .full
		.empty       (empty),       //            .empty
		.almost_full (almost_full)  //            .almost_full
	);

endmodule
