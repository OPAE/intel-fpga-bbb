// mult_8bit.v

// Generated using ACDS version 16.0 211

`timescale 1 ps / 1 ps
module mult_8bit (
		input  wire [7:0]  dataa,  //  mult_input.dataa
		input  wire [7:0]  datab,  //            .datab
		input  wire        clock,  //            .clock
        input  wire        clken,  //            .clken
		input  wire        aclr,   //            .aclr
		output wire [15:0] result  // mult_output.result
	);

	mult_8bit_lpm_mult_160_lkaps7i lpm_mult_0 (
		.dataa  (dataa),  //  mult_input.dataa
		.datab  (datab),  //            .datab
		.clock  (clock),  //            .clock
        .clken  (clken),  //            .clken
		.aclr   (aclr),   //            .aclr
		.result (result)  // mult_output.result
	);

endmodule
